module Adder(
  input         io_cin,
  input  [31:0] io_A_in,
  input  [31:0] io_B_in,
  output        io_zero,
  output        io_carry,
  output        io_overflow,
  output        io_negative,
  output [31:0] io_O_out
);
  wire [31:0] _B_in_not_T_1 = ~io_B_in; // @[Adder.scala 19:38]
  wire [31:0] B_in_not = io_cin ? _B_in_not_T_1 : io_B_in; // @[Adder.scala 19:23]
  wire [32:0] _res_T = io_A_in + B_in_not; // @[Adder.scala 20:23]
  wire [32:0] _GEN_0 = {{32'd0}, io_cin}; // @[Adder.scala 20:35]
  wire [33:0] res = _res_T + _GEN_0; // @[Adder.scala 20:35]
  assign io_zero = io_O_out == 32'h0; // @[Adder.scala 26:26]
  assign io_carry = res[32]; // @[Adder.scala 22:20]
  assign io_overflow = io_A_in[31] & B_in_not[31] & ~res[31] | ~io_A_in[31] & ~B_in_not[31] & res[31]; // @[Adder.scala 24:62]
  assign io_negative = res[31]; // @[Adder.scala 25:23]
  assign io_O_out = res[31:0]; // @[Adder.scala 23:20]
endmodule
module ALU(
  input         clock,
  input         reset,
  input  [31:0] io_A_in,
  input  [31:0] io_B_in,
  input  [3:0]  io_ALU_op,
  output [31:0] io_ALU_out,
  output        io_Zero,
  output        io_Less,
  output        io_Overflow_out
);
  wire  adder_io_cin; // @[ALU.scala 26:23]
  wire [31:0] adder_io_A_in; // @[ALU.scala 26:23]
  wire [31:0] adder_io_B_in; // @[ALU.scala 26:23]
  wire  adder_io_zero; // @[ALU.scala 26:23]
  wire  adder_io_carry; // @[ALU.scala 26:23]
  wire  adder_io_overflow; // @[ALU.scala 26:23]
  wire  adder_io_negative; // @[ALU.scala 26:23]
  wire [31:0] adder_io_O_out; // @[ALU.scala 26:23]
  wire  _ctrl_T_1 = ~io_ALU_op[3]; // @[ALU.scala 19:10]
  wire  _ctrl_T_3 = ~io_ALU_op[1]; // @[ALU.scala 19:26]
  wire  _ctrl_T_10 = ~io_ALU_op[3] & io_ALU_op[2] & io_ALU_op[0]; // @[ALU.scala 19:73]
  wire  _ctrl_T_14 = io_ALU_op[3] & io_ALU_op[1]; // @[ALU.scala 19:105]
  wire  ctrl_hi = ~io_ALU_op[3] & ~io_ALU_op[1] | ~io_ALU_op[3] & io_ALU_op[2] & io_ALU_op[0] | io_ALU_op[3] & io_ALU_op
    [1]; // @[ALU.scala 19:89]
  wire  _ctrl_T_18 = ~io_ALU_op[2]; // @[ALU.scala 21:30]
  wire  ctrl_hi_1 = _ctrl_T_1 & ~io_ALU_op[2] & _ctrl_T_3 | io_ALU_op[3] & ~io_ALU_op[2] & ~io_ALU_op[0] | io_ALU_op[2]
     & io_ALU_op[1] & ~io_ALU_op[0] | _ctrl_T_14; // @[ALU.scala 21:158]
  wire  ctrl_lo = _ctrl_T_18 & _ctrl_T_3 | _ctrl_T_10 | io_ALU_op[3] & io_ALU_op[2] & io_ALU_op[1]; // @[ALU.scala 22:93]
  wire [2:0] ctrl = {ctrl_hi,ctrl_hi_1,ctrl_lo}; // @[Cat.scala 30:58]
  wire [31:0] _A_in_not_T_1 = ~io_A_in; // @[ALU.scala 44:38]
  wire [31:0] A_in_not = io_ALU_op[0] ? _A_in_not_T_1 : io_A_in; // @[ALU.scala 44:23]
  wire  tocount_31 = ~A_in_not[31]; // @[ALU.scala 48:45]
  wire  tocount_30 = tocount_31 & ~A_in_not[30]; // @[ALU.scala 49:41]
  wire  tocount_29 = tocount_30 & ~A_in_not[29]; // @[ALU.scala 49:41]
  wire  tocount_28 = tocount_29 & ~A_in_not[28]; // @[ALU.scala 49:41]
  wire  tocount_27 = tocount_28 & ~A_in_not[27]; // @[ALU.scala 49:41]
  wire  tocount_26 = tocount_27 & ~A_in_not[26]; // @[ALU.scala 49:41]
  wire  tocount_25 = tocount_26 & ~A_in_not[25]; // @[ALU.scala 49:41]
  wire  tocount_24 = tocount_25 & ~A_in_not[24]; // @[ALU.scala 49:41]
  wire  tocount_23 = tocount_24 & ~A_in_not[23]; // @[ALU.scala 49:41]
  wire  tocount_22 = tocount_23 & ~A_in_not[22]; // @[ALU.scala 49:41]
  wire  tocount_21 = tocount_22 & ~A_in_not[21]; // @[ALU.scala 49:41]
  wire  tocount_20 = tocount_21 & ~A_in_not[20]; // @[ALU.scala 49:41]
  wire  tocount_19 = tocount_20 & ~A_in_not[19]; // @[ALU.scala 49:41]
  wire  tocount_18 = tocount_19 & ~A_in_not[18]; // @[ALU.scala 49:41]
  wire  tocount_17 = tocount_18 & ~A_in_not[17]; // @[ALU.scala 49:41]
  wire  tocount_16 = tocount_17 & ~A_in_not[16]; // @[ALU.scala 49:41]
  wire  tocount_15 = tocount_16 & ~A_in_not[15]; // @[ALU.scala 49:41]
  wire  tocount_14 = tocount_15 & ~A_in_not[14]; // @[ALU.scala 49:41]
  wire  tocount_13 = tocount_14 & ~A_in_not[13]; // @[ALU.scala 49:41]
  wire  tocount_12 = tocount_13 & ~A_in_not[12]; // @[ALU.scala 49:41]
  wire  tocount_11 = tocount_12 & ~A_in_not[11]; // @[ALU.scala 49:41]
  wire  tocount_10 = tocount_11 & ~A_in_not[10]; // @[ALU.scala 49:41]
  wire  tocount_9 = tocount_10 & ~A_in_not[9]; // @[ALU.scala 49:41]
  wire  tocount_8 = tocount_9 & ~A_in_not[8]; // @[ALU.scala 49:41]
  wire  tocount_7 = tocount_8 & ~A_in_not[7]; // @[ALU.scala 49:41]
  wire  tocount_6 = tocount_7 & ~A_in_not[6]; // @[ALU.scala 49:41]
  wire  tocount_5 = tocount_6 & ~A_in_not[5]; // @[ALU.scala 49:41]
  wire  tocount_4 = tocount_5 & ~A_in_not[4]; // @[ALU.scala 49:41]
  wire  tocount_3 = tocount_4 & ~A_in_not[3]; // @[ALU.scala 49:41]
  wire  tocount_2 = tocount_3 & ~A_in_not[2]; // @[ALU.scala 49:41]
  wire  tocount_1 = tocount_2 & ~A_in_not[1]; // @[ALU.scala 49:41]
  wire  tocount_0 = tocount_1 & ~A_in_not[0]; // @[ALU.scala 49:41]
  wire [5:0] count_31 = {{5'd0}, tocount_31}; // @[ALU.scala 46:21 ALU.scala 52:28]
  wire [5:0] _count_30_T_1 = count_31 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_30 = tocount_30 ? _count_30_T_1 : count_31; // @[ALU.scala 53:29]
  wire [5:0] _count_29_T_1 = count_30 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_29 = tocount_29 ? _count_29_T_1 : count_30; // @[ALU.scala 53:29]
  wire [5:0] _count_28_T_1 = count_29 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_28 = tocount_28 ? _count_28_T_1 : count_29; // @[ALU.scala 53:29]
  wire [5:0] _count_27_T_1 = count_28 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_27 = tocount_27 ? _count_27_T_1 : count_28; // @[ALU.scala 53:29]
  wire [5:0] _count_26_T_1 = count_27 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_26 = tocount_26 ? _count_26_T_1 : count_27; // @[ALU.scala 53:29]
  wire [5:0] _count_25_T_1 = count_26 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_25 = tocount_25 ? _count_25_T_1 : count_26; // @[ALU.scala 53:29]
  wire [5:0] _count_24_T_1 = count_25 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_24 = tocount_24 ? _count_24_T_1 : count_25; // @[ALU.scala 53:29]
  wire [5:0] _count_23_T_1 = count_24 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_23 = tocount_23 ? _count_23_T_1 : count_24; // @[ALU.scala 53:29]
  wire [5:0] _count_22_T_1 = count_23 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_22 = tocount_22 ? _count_22_T_1 : count_23; // @[ALU.scala 53:29]
  wire [5:0] _count_21_T_1 = count_22 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_21 = tocount_21 ? _count_21_T_1 : count_22; // @[ALU.scala 53:29]
  wire [5:0] _count_20_T_1 = count_21 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_20 = tocount_20 ? _count_20_T_1 : count_21; // @[ALU.scala 53:29]
  wire [5:0] _count_19_T_1 = count_20 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_19 = tocount_19 ? _count_19_T_1 : count_20; // @[ALU.scala 53:29]
  wire [5:0] _count_18_T_1 = count_19 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_18 = tocount_18 ? _count_18_T_1 : count_19; // @[ALU.scala 53:29]
  wire [5:0] _count_17_T_1 = count_18 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_17 = tocount_17 ? _count_17_T_1 : count_18; // @[ALU.scala 53:29]
  wire [5:0] _count_16_T_1 = count_17 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_16 = tocount_16 ? _count_16_T_1 : count_17; // @[ALU.scala 53:29]
  wire [5:0] _count_15_T_1 = count_16 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_15 = tocount_15 ? _count_15_T_1 : count_16; // @[ALU.scala 53:29]
  wire [5:0] _count_14_T_1 = count_15 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_14 = tocount_14 ? _count_14_T_1 : count_15; // @[ALU.scala 53:29]
  wire [5:0] _count_13_T_1 = count_14 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_13 = tocount_13 ? _count_13_T_1 : count_14; // @[ALU.scala 53:29]
  wire [5:0] _count_12_T_1 = count_13 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_12 = tocount_12 ? _count_12_T_1 : count_13; // @[ALU.scala 53:29]
  wire [5:0] _count_11_T_1 = count_12 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_11 = tocount_11 ? _count_11_T_1 : count_12; // @[ALU.scala 53:29]
  wire [5:0] _count_10_T_1 = count_11 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_10 = tocount_10 ? _count_10_T_1 : count_11; // @[ALU.scala 53:29]
  wire [5:0] _count_9_T_1 = count_10 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_9 = tocount_9 ? _count_9_T_1 : count_10; // @[ALU.scala 53:29]
  wire [5:0] _count_8_T_1 = count_9 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_8 = tocount_8 ? _count_8_T_1 : count_9; // @[ALU.scala 53:29]
  wire [5:0] _count_7_T_1 = count_8 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_7 = tocount_7 ? _count_7_T_1 : count_8; // @[ALU.scala 53:29]
  wire [5:0] _count_6_T_1 = count_7 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_6 = tocount_6 ? _count_6_T_1 : count_7; // @[ALU.scala 53:29]
  wire [5:0] _count_5_T_1 = count_6 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_5 = tocount_5 ? _count_5_T_1 : count_6; // @[ALU.scala 53:29]
  wire [5:0] _count_4_T_1 = count_5 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_4 = tocount_4 ? _count_4_T_1 : count_5; // @[ALU.scala 53:29]
  wire [5:0] _count_3_T_1 = count_4 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_3 = tocount_3 ? _count_3_T_1 : count_4; // @[ALU.scala 53:29]
  wire [5:0] _count_2_T_1 = count_3 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_2 = tocount_2 ? _count_2_T_1 : count_3; // @[ALU.scala 53:29]
  wire [5:0] _count_1_T_1 = count_2 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_1 = tocount_1 ? _count_1_T_1 : count_2; // @[ALU.scala 53:29]
  wire [5:0] _count_0_T_1 = count_1 + 6'h1; // @[ALU.scala 53:52]
  wire [5:0] count_0 = tocount_0 ? _count_0_T_1 : count_1; // @[ALU.scala 53:29]
  wire [31:0] _io_ALU_out_T = io_A_in ^ io_B_in; // @[ALU.scala 60:31]
  wire [31:0] _io_ALU_out_T_1 = io_A_in | io_B_in; // @[ALU.scala 62:31]
  wire [31:0] _io_ALU_out_T_3 = ~_io_ALU_out_T_1; // @[ALU.scala 64:23]
  wire [31:0] _io_ALU_out_T_4 = io_A_in & io_B_in; // @[ALU.scala 66:31]
  wire [15:0] io_ALU_out_hi = io_B_in[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] io_ALU_out_lo = io_B_in[15:0]; // @[ALU.scala 71:51]
  wire [31:0] _io_ALU_out_T_9 = {io_ALU_out_hi,io_ALU_out_lo}; // @[Cat.scala 30:58]
  wire [23:0] io_ALU_out_hi_1 = io_B_in[7] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_ALU_out_lo_1 = io_B_in[7:0]; // @[ALU.scala 72:50]
  wire [31:0] _io_ALU_out_T_12 = {io_ALU_out_hi_1,io_ALU_out_lo_1}; // @[Cat.scala 30:58]
  wire [31:0] _io_ALU_out_T_13 = io_ALU_op[0] ? _io_ALU_out_T_9 : _io_ALU_out_T_12; // @[ALU.scala 70:26]
  wire [31:0] _GEN_2 = ctrl == 3'h7 ? adder_io_O_out : 32'h0; // @[ALU.scala 74:32 ALU.scala 75:20 ALU.scala 56:16]
  wire [31:0] _GEN_3 = ctrl == 3'h6 ? _io_ALU_out_T_13 : _GEN_2; // @[ALU.scala 69:31 ALU.scala 70:20]
  wire [31:0] _GEN_4 = ctrl == 3'h5 ? {{31'd0}, io_Less} : _GEN_3; // @[ALU.scala 67:31 ALU.scala 68:20]
  wire [31:0] _GEN_5 = ctrl == 3'h4 ? _io_ALU_out_T_4 : _GEN_4; // @[ALU.scala 65:32 ALU.scala 66:20]
  wire [31:0] _GEN_6 = ctrl == 3'h3 ? _io_ALU_out_T_3 : _GEN_5; // @[ALU.scala 63:31 ALU.scala 64:20]
  wire [31:0] _GEN_7 = ctrl == 3'h2 ? _io_ALU_out_T_1 : _GEN_6; // @[ALU.scala 61:32 ALU.scala 62:20]
  wire [31:0] _GEN_8 = ctrl == 3'h1 ? _io_ALU_out_T : _GEN_7; // @[ALU.scala 59:30 ALU.scala 60:20]
  Adder adder ( // @[ALU.scala 26:23]
    .io_cin(adder_io_cin),
    .io_A_in(adder_io_A_in),
    .io_B_in(adder_io_B_in),
    .io_zero(adder_io_zero),
    .io_carry(adder_io_carry),
    .io_overflow(adder_io_overflow),
    .io_negative(adder_io_negative),
    .io_O_out(adder_io_O_out)
  );
  assign io_ALU_out = ctrl == 3'h0 ? {{26'd0}, count_0} : _GEN_8; // @[ALU.scala 57:24 ALU.scala 58:20]
  assign io_Zero = adder_io_zero; // @[ALU.scala 30:13]
  assign io_Less = io_ALU_op == 4'h7 ? ~adder_io_carry : adder_io_overflow ^ adder_io_negative; // @[ALU.scala 38:26 ALU.scala 39:17 ALU.scala 41:17]
  assign io_Overflow_out = io_ALU_op[3:1] == 3'h7 & adder_io_overflow; // @[ALU.scala 32:34 ALU.scala 33:25 ALU.scala 35:25]
  assign adder_io_cin = io_ALU_op[0]; // @[ALU.scala 29:30]
  assign adder_io_A_in = io_A_in; // @[ALU.scala 27:19]
  assign adder_io_B_in = io_B_in; // @[ALU.scala 28:19]
endmodule

module Register(
  input         clock,
  input         reset,
  input  [4:0]  io_Rs_addr,
  input  [4:0]  io_Rt_addr,
  input  [4:0]  io_Rd_addr,
  input  [31:0] io_Rd_in,
  input  [3:0]  io_Rd_byte_w_en,
  output [31:0] io_Rs_out,
  output [31:0] io_Rt_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] reg_0_0; // @[Register.scala 17:22]
  reg [7:0] reg_0_1; // @[Register.scala 17:22]
  reg [7:0] reg_0_2; // @[Register.scala 17:22]
  reg [7:0] reg_0_3; // @[Register.scala 17:22]
  reg [7:0] reg_1_0; // @[Register.scala 17:22]
  reg [7:0] reg_1_1; // @[Register.scala 17:22]
  reg [7:0] reg_1_2; // @[Register.scala 17:22]
  reg [7:0] reg_1_3; // @[Register.scala 17:22]
  reg [7:0] reg_2_0; // @[Register.scala 17:22]
  reg [7:0] reg_2_1; // @[Register.scala 17:22]
  reg [7:0] reg_2_2; // @[Register.scala 17:22]
  reg [7:0] reg_2_3; // @[Register.scala 17:22]
  reg [7:0] reg_3_0; // @[Register.scala 17:22]
  reg [7:0] reg_3_1; // @[Register.scala 17:22]
  reg [7:0] reg_3_2; // @[Register.scala 17:22]
  reg [7:0] reg_3_3; // @[Register.scala 17:22]
  reg [7:0] reg_4_0; // @[Register.scala 17:22]
  reg [7:0] reg_4_1; // @[Register.scala 17:22]
  reg [7:0] reg_4_2; // @[Register.scala 17:22]
  reg [7:0] reg_4_3; // @[Register.scala 17:22]
  reg [7:0] reg_5_0; // @[Register.scala 17:22]
  reg [7:0] reg_5_1; // @[Register.scala 17:22]
  reg [7:0] reg_5_2; // @[Register.scala 17:22]
  reg [7:0] reg_5_3; // @[Register.scala 17:22]
  reg [7:0] reg_6_0; // @[Register.scala 17:22]
  reg [7:0] reg_6_1; // @[Register.scala 17:22]
  reg [7:0] reg_6_2; // @[Register.scala 17:22]
  reg [7:0] reg_6_3; // @[Register.scala 17:22]
  reg [7:0] reg_7_0; // @[Register.scala 17:22]
  reg [7:0] reg_7_1; // @[Register.scala 17:22]
  reg [7:0] reg_7_2; // @[Register.scala 17:22]
  reg [7:0] reg_7_3; // @[Register.scala 17:22]
  reg [7:0] reg_8_0; // @[Register.scala 17:22]
  reg [7:0] reg_8_1; // @[Register.scala 17:22]
  reg [7:0] reg_8_2; // @[Register.scala 17:22]
  reg [7:0] reg_8_3; // @[Register.scala 17:22]
  reg [7:0] reg_9_0; // @[Register.scala 17:22]
  reg [7:0] reg_9_1; // @[Register.scala 17:22]
  reg [7:0] reg_9_2; // @[Register.scala 17:22]
  reg [7:0] reg_9_3; // @[Register.scala 17:22]
  reg [7:0] reg_10_0; // @[Register.scala 17:22]
  reg [7:0] reg_10_1; // @[Register.scala 17:22]
  reg [7:0] reg_10_2; // @[Register.scala 17:22]
  reg [7:0] reg_10_3; // @[Register.scala 17:22]
  reg [7:0] reg_11_0; // @[Register.scala 17:22]
  reg [7:0] reg_11_1; // @[Register.scala 17:22]
  reg [7:0] reg_11_2; // @[Register.scala 17:22]
  reg [7:0] reg_11_3; // @[Register.scala 17:22]
  reg [7:0] reg_12_0; // @[Register.scala 17:22]
  reg [7:0] reg_12_1; // @[Register.scala 17:22]
  reg [7:0] reg_12_2; // @[Register.scala 17:22]
  reg [7:0] reg_12_3; // @[Register.scala 17:22]
  reg [7:0] reg_13_0; // @[Register.scala 17:22]
  reg [7:0] reg_13_1; // @[Register.scala 17:22]
  reg [7:0] reg_13_2; // @[Register.scala 17:22]
  reg [7:0] reg_13_3; // @[Register.scala 17:22]
  reg [7:0] reg_14_0; // @[Register.scala 17:22]
  reg [7:0] reg_14_1; // @[Register.scala 17:22]
  reg [7:0] reg_14_2; // @[Register.scala 17:22]
  reg [7:0] reg_14_3; // @[Register.scala 17:22]
  reg [7:0] reg_15_0; // @[Register.scala 17:22]
  reg [7:0] reg_15_1; // @[Register.scala 17:22]
  reg [7:0] reg_15_2; // @[Register.scala 17:22]
  reg [7:0] reg_15_3; // @[Register.scala 17:22]
  reg [7:0] reg_16_0; // @[Register.scala 17:22]
  reg [7:0] reg_16_1; // @[Register.scala 17:22]
  reg [7:0] reg_16_2; // @[Register.scala 17:22]
  reg [7:0] reg_16_3; // @[Register.scala 17:22]
  reg [7:0] reg_17_0; // @[Register.scala 17:22]
  reg [7:0] reg_17_1; // @[Register.scala 17:22]
  reg [7:0] reg_17_2; // @[Register.scala 17:22]
  reg [7:0] reg_17_3; // @[Register.scala 17:22]
  reg [7:0] reg_18_0; // @[Register.scala 17:22]
  reg [7:0] reg_18_1; // @[Register.scala 17:22]
  reg [7:0] reg_18_2; // @[Register.scala 17:22]
  reg [7:0] reg_18_3; // @[Register.scala 17:22]
  reg [7:0] reg_19_0; // @[Register.scala 17:22]
  reg [7:0] reg_19_1; // @[Register.scala 17:22]
  reg [7:0] reg_19_2; // @[Register.scala 17:22]
  reg [7:0] reg_19_3; // @[Register.scala 17:22]
  reg [7:0] reg_20_0; // @[Register.scala 17:22]
  reg [7:0] reg_20_1; // @[Register.scala 17:22]
  reg [7:0] reg_20_2; // @[Register.scala 17:22]
  reg [7:0] reg_20_3; // @[Register.scala 17:22]
  reg [7:0] reg_21_0; // @[Register.scala 17:22]
  reg [7:0] reg_21_1; // @[Register.scala 17:22]
  reg [7:0] reg_21_2; // @[Register.scala 17:22]
  reg [7:0] reg_21_3; // @[Register.scala 17:22]
  reg [7:0] reg_22_0; // @[Register.scala 17:22]
  reg [7:0] reg_22_1; // @[Register.scala 17:22]
  reg [7:0] reg_22_2; // @[Register.scala 17:22]
  reg [7:0] reg_22_3; // @[Register.scala 17:22]
  reg [7:0] reg_23_0; // @[Register.scala 17:22]
  reg [7:0] reg_23_1; // @[Register.scala 17:22]
  reg [7:0] reg_23_2; // @[Register.scala 17:22]
  reg [7:0] reg_23_3; // @[Register.scala 17:22]
  reg [7:0] reg_24_0; // @[Register.scala 17:22]
  reg [7:0] reg_24_1; // @[Register.scala 17:22]
  reg [7:0] reg_24_2; // @[Register.scala 17:22]
  reg [7:0] reg_24_3; // @[Register.scala 17:22]
  reg [7:0] reg_25_0; // @[Register.scala 17:22]
  reg [7:0] reg_25_1; // @[Register.scala 17:22]
  reg [7:0] reg_25_2; // @[Register.scala 17:22]
  reg [7:0] reg_25_3; // @[Register.scala 17:22]
  reg [7:0] reg_26_0; // @[Register.scala 17:22]
  reg [7:0] reg_26_1; // @[Register.scala 17:22]
  reg [7:0] reg_26_2; // @[Register.scala 17:22]
  reg [7:0] reg_26_3; // @[Register.scala 17:22]
  reg [7:0] reg_27_0; // @[Register.scala 17:22]
  reg [7:0] reg_27_1; // @[Register.scala 17:22]
  reg [7:0] reg_27_2; // @[Register.scala 17:22]
  reg [7:0] reg_27_3; // @[Register.scala 17:22]
  reg [7:0] reg_28_0; // @[Register.scala 17:22]
  reg [7:0] reg_28_1; // @[Register.scala 17:22]
  reg [7:0] reg_28_2; // @[Register.scala 17:22]
  reg [7:0] reg_28_3; // @[Register.scala 17:22]
  reg [7:0] reg_29_0; // @[Register.scala 17:22]
  reg [7:0] reg_29_1; // @[Register.scala 17:22]
  reg [7:0] reg_29_2; // @[Register.scala 17:22]
  reg [7:0] reg_29_3; // @[Register.scala 17:22]
  reg [7:0] reg_30_0; // @[Register.scala 17:22]
  reg [7:0] reg_30_1; // @[Register.scala 17:22]
  reg [7:0] reg_30_2; // @[Register.scala 17:22]
  reg [7:0] reg_30_3; // @[Register.scala 17:22]
  reg [7:0] reg_31_0; // @[Register.scala 17:22]
  reg [7:0] reg_31_1; // @[Register.scala 17:22]
  reg [7:0] reg_31_2; // @[Register.scala 17:22]
  reg [7:0] reg_31_3; // @[Register.scala 17:22]
  wire [7:0] _GEN_1 = 5'h1 == io_Rs_addr ? reg_1_3 : reg_0_3; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_2 = 5'h2 == io_Rs_addr ? reg_2_3 : _GEN_1; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_3 = 5'h3 == io_Rs_addr ? reg_3_3 : _GEN_2; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_4 = 5'h4 == io_Rs_addr ? reg_4_3 : _GEN_3; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_5 = 5'h5 == io_Rs_addr ? reg_5_3 : _GEN_4; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_6 = 5'h6 == io_Rs_addr ? reg_6_3 : _GEN_5; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_7 = 5'h7 == io_Rs_addr ? reg_7_3 : _GEN_6; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_8 = 5'h8 == io_Rs_addr ? reg_8_3 : _GEN_7; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_9 = 5'h9 == io_Rs_addr ? reg_9_3 : _GEN_8; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_10 = 5'ha == io_Rs_addr ? reg_10_3 : _GEN_9; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_11 = 5'hb == io_Rs_addr ? reg_11_3 : _GEN_10; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_12 = 5'hc == io_Rs_addr ? reg_12_3 : _GEN_11; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_13 = 5'hd == io_Rs_addr ? reg_13_3 : _GEN_12; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_14 = 5'he == io_Rs_addr ? reg_14_3 : _GEN_13; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_15 = 5'hf == io_Rs_addr ? reg_15_3 : _GEN_14; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_16 = 5'h10 == io_Rs_addr ? reg_16_3 : _GEN_15; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_17 = 5'h11 == io_Rs_addr ? reg_17_3 : _GEN_16; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_18 = 5'h12 == io_Rs_addr ? reg_18_3 : _GEN_17; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_19 = 5'h13 == io_Rs_addr ? reg_19_3 : _GEN_18; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_20 = 5'h14 == io_Rs_addr ? reg_20_3 : _GEN_19; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_21 = 5'h15 == io_Rs_addr ? reg_21_3 : _GEN_20; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_22 = 5'h16 == io_Rs_addr ? reg_22_3 : _GEN_21; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_23 = 5'h17 == io_Rs_addr ? reg_23_3 : _GEN_22; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_24 = 5'h18 == io_Rs_addr ? reg_24_3 : _GEN_23; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_25 = 5'h19 == io_Rs_addr ? reg_25_3 : _GEN_24; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_26 = 5'h1a == io_Rs_addr ? reg_26_3 : _GEN_25; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_27 = 5'h1b == io_Rs_addr ? reg_27_3 : _GEN_26; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_28 = 5'h1c == io_Rs_addr ? reg_28_3 : _GEN_27; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_29 = 5'h1d == io_Rs_addr ? reg_29_3 : _GEN_28; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_30 = 5'h1e == io_Rs_addr ? reg_30_3 : _GEN_29; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_31 = 5'h1f == io_Rs_addr ? reg_31_3 : _GEN_30; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_33 = 5'h1 == io_Rs_addr ? reg_1_2 : reg_0_2; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_34 = 5'h2 == io_Rs_addr ? reg_2_2 : _GEN_33; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_35 = 5'h3 == io_Rs_addr ? reg_3_2 : _GEN_34; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_36 = 5'h4 == io_Rs_addr ? reg_4_2 : _GEN_35; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_37 = 5'h5 == io_Rs_addr ? reg_5_2 : _GEN_36; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_38 = 5'h6 == io_Rs_addr ? reg_6_2 : _GEN_37; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_39 = 5'h7 == io_Rs_addr ? reg_7_2 : _GEN_38; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_40 = 5'h8 == io_Rs_addr ? reg_8_2 : _GEN_39; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_41 = 5'h9 == io_Rs_addr ? reg_9_2 : _GEN_40; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_42 = 5'ha == io_Rs_addr ? reg_10_2 : _GEN_41; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_43 = 5'hb == io_Rs_addr ? reg_11_2 : _GEN_42; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_44 = 5'hc == io_Rs_addr ? reg_12_2 : _GEN_43; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_45 = 5'hd == io_Rs_addr ? reg_13_2 : _GEN_44; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_46 = 5'he == io_Rs_addr ? reg_14_2 : _GEN_45; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_47 = 5'hf == io_Rs_addr ? reg_15_2 : _GEN_46; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_48 = 5'h10 == io_Rs_addr ? reg_16_2 : _GEN_47; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_49 = 5'h11 == io_Rs_addr ? reg_17_2 : _GEN_48; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_50 = 5'h12 == io_Rs_addr ? reg_18_2 : _GEN_49; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_51 = 5'h13 == io_Rs_addr ? reg_19_2 : _GEN_50; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_52 = 5'h14 == io_Rs_addr ? reg_20_2 : _GEN_51; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_53 = 5'h15 == io_Rs_addr ? reg_21_2 : _GEN_52; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_54 = 5'h16 == io_Rs_addr ? reg_22_2 : _GEN_53; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_55 = 5'h17 == io_Rs_addr ? reg_23_2 : _GEN_54; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_56 = 5'h18 == io_Rs_addr ? reg_24_2 : _GEN_55; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_57 = 5'h19 == io_Rs_addr ? reg_25_2 : _GEN_56; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_58 = 5'h1a == io_Rs_addr ? reg_26_2 : _GEN_57; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_59 = 5'h1b == io_Rs_addr ? reg_27_2 : _GEN_58; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_60 = 5'h1c == io_Rs_addr ? reg_28_2 : _GEN_59; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_61 = 5'h1d == io_Rs_addr ? reg_29_2 : _GEN_60; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_62 = 5'h1e == io_Rs_addr ? reg_30_2 : _GEN_61; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_63 = 5'h1f == io_Rs_addr ? reg_31_2 : _GEN_62; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_65 = 5'h1 == io_Rs_addr ? reg_1_1 : reg_0_1; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_66 = 5'h2 == io_Rs_addr ? reg_2_1 : _GEN_65; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_67 = 5'h3 == io_Rs_addr ? reg_3_1 : _GEN_66; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_68 = 5'h4 == io_Rs_addr ? reg_4_1 : _GEN_67; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_69 = 5'h5 == io_Rs_addr ? reg_5_1 : _GEN_68; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_70 = 5'h6 == io_Rs_addr ? reg_6_1 : _GEN_69; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_71 = 5'h7 == io_Rs_addr ? reg_7_1 : _GEN_70; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_72 = 5'h8 == io_Rs_addr ? reg_8_1 : _GEN_71; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_73 = 5'h9 == io_Rs_addr ? reg_9_1 : _GEN_72; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_74 = 5'ha == io_Rs_addr ? reg_10_1 : _GEN_73; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_75 = 5'hb == io_Rs_addr ? reg_11_1 : _GEN_74; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_76 = 5'hc == io_Rs_addr ? reg_12_1 : _GEN_75; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_77 = 5'hd == io_Rs_addr ? reg_13_1 : _GEN_76; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_78 = 5'he == io_Rs_addr ? reg_14_1 : _GEN_77; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_79 = 5'hf == io_Rs_addr ? reg_15_1 : _GEN_78; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_80 = 5'h10 == io_Rs_addr ? reg_16_1 : _GEN_79; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_81 = 5'h11 == io_Rs_addr ? reg_17_1 : _GEN_80; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_82 = 5'h12 == io_Rs_addr ? reg_18_1 : _GEN_81; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_83 = 5'h13 == io_Rs_addr ? reg_19_1 : _GEN_82; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_84 = 5'h14 == io_Rs_addr ? reg_20_1 : _GEN_83; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_85 = 5'h15 == io_Rs_addr ? reg_21_1 : _GEN_84; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_86 = 5'h16 == io_Rs_addr ? reg_22_1 : _GEN_85; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_87 = 5'h17 == io_Rs_addr ? reg_23_1 : _GEN_86; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_88 = 5'h18 == io_Rs_addr ? reg_24_1 : _GEN_87; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_89 = 5'h19 == io_Rs_addr ? reg_25_1 : _GEN_88; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_90 = 5'h1a == io_Rs_addr ? reg_26_1 : _GEN_89; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_91 = 5'h1b == io_Rs_addr ? reg_27_1 : _GEN_90; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_92 = 5'h1c == io_Rs_addr ? reg_28_1 : _GEN_91; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_93 = 5'h1d == io_Rs_addr ? reg_29_1 : _GEN_92; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_94 = 5'h1e == io_Rs_addr ? reg_30_1 : _GEN_93; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_95 = 5'h1f == io_Rs_addr ? reg_31_1 : _GEN_94; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [23:0] io_Rs_out_hi_1 = {_GEN_31,_GEN_63,_GEN_95}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_97 = 5'h1 == io_Rs_addr ? reg_1_0 : reg_0_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_98 = 5'h2 == io_Rs_addr ? reg_2_0 : _GEN_97; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_99 = 5'h3 == io_Rs_addr ? reg_3_0 : _GEN_98; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_100 = 5'h4 == io_Rs_addr ? reg_4_0 : _GEN_99; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_101 = 5'h5 == io_Rs_addr ? reg_5_0 : _GEN_100; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_102 = 5'h6 == io_Rs_addr ? reg_6_0 : _GEN_101; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_103 = 5'h7 == io_Rs_addr ? reg_7_0 : _GEN_102; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_104 = 5'h8 == io_Rs_addr ? reg_8_0 : _GEN_103; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_105 = 5'h9 == io_Rs_addr ? reg_9_0 : _GEN_104; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_106 = 5'ha == io_Rs_addr ? reg_10_0 : _GEN_105; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_107 = 5'hb == io_Rs_addr ? reg_11_0 : _GEN_106; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_108 = 5'hc == io_Rs_addr ? reg_12_0 : _GEN_107; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_109 = 5'hd == io_Rs_addr ? reg_13_0 : _GEN_108; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_110 = 5'he == io_Rs_addr ? reg_14_0 : _GEN_109; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_111 = 5'hf == io_Rs_addr ? reg_15_0 : _GEN_110; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_112 = 5'h10 == io_Rs_addr ? reg_16_0 : _GEN_111; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_113 = 5'h11 == io_Rs_addr ? reg_17_0 : _GEN_112; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_114 = 5'h12 == io_Rs_addr ? reg_18_0 : _GEN_113; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_115 = 5'h13 == io_Rs_addr ? reg_19_0 : _GEN_114; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_116 = 5'h14 == io_Rs_addr ? reg_20_0 : _GEN_115; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_117 = 5'h15 == io_Rs_addr ? reg_21_0 : _GEN_116; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_118 = 5'h16 == io_Rs_addr ? reg_22_0 : _GEN_117; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_119 = 5'h17 == io_Rs_addr ? reg_23_0 : _GEN_118; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_120 = 5'h18 == io_Rs_addr ? reg_24_0 : _GEN_119; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_121 = 5'h19 == io_Rs_addr ? reg_25_0 : _GEN_120; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_122 = 5'h1a == io_Rs_addr ? reg_26_0 : _GEN_121; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_123 = 5'h1b == io_Rs_addr ? reg_27_0 : _GEN_122; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_124 = 5'h1c == io_Rs_addr ? reg_28_0 : _GEN_123; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_125 = 5'h1d == io_Rs_addr ? reg_29_0 : _GEN_124; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_126 = 5'h1e == io_Rs_addr ? reg_30_0 : _GEN_125; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_127 = 5'h1f == io_Rs_addr ? reg_31_0 : _GEN_126; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_129 = 5'h1 == io_Rt_addr ? reg_1_3 : reg_0_3; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_130 = 5'h2 == io_Rt_addr ? reg_2_3 : _GEN_129; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_131 = 5'h3 == io_Rt_addr ? reg_3_3 : _GEN_130; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_132 = 5'h4 == io_Rt_addr ? reg_4_3 : _GEN_131; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_133 = 5'h5 == io_Rt_addr ? reg_5_3 : _GEN_132; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_134 = 5'h6 == io_Rt_addr ? reg_6_3 : _GEN_133; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_135 = 5'h7 == io_Rt_addr ? reg_7_3 : _GEN_134; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_136 = 5'h8 == io_Rt_addr ? reg_8_3 : _GEN_135; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_137 = 5'h9 == io_Rt_addr ? reg_9_3 : _GEN_136; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_138 = 5'ha == io_Rt_addr ? reg_10_3 : _GEN_137; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_139 = 5'hb == io_Rt_addr ? reg_11_3 : _GEN_138; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_140 = 5'hc == io_Rt_addr ? reg_12_3 : _GEN_139; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_141 = 5'hd == io_Rt_addr ? reg_13_3 : _GEN_140; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_142 = 5'he == io_Rt_addr ? reg_14_3 : _GEN_141; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_143 = 5'hf == io_Rt_addr ? reg_15_3 : _GEN_142; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_144 = 5'h10 == io_Rt_addr ? reg_16_3 : _GEN_143; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_145 = 5'h11 == io_Rt_addr ? reg_17_3 : _GEN_144; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_146 = 5'h12 == io_Rt_addr ? reg_18_3 : _GEN_145; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_147 = 5'h13 == io_Rt_addr ? reg_19_3 : _GEN_146; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_148 = 5'h14 == io_Rt_addr ? reg_20_3 : _GEN_147; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_149 = 5'h15 == io_Rt_addr ? reg_21_3 : _GEN_148; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_150 = 5'h16 == io_Rt_addr ? reg_22_3 : _GEN_149; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_151 = 5'h17 == io_Rt_addr ? reg_23_3 : _GEN_150; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_152 = 5'h18 == io_Rt_addr ? reg_24_3 : _GEN_151; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_153 = 5'h19 == io_Rt_addr ? reg_25_3 : _GEN_152; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_154 = 5'h1a == io_Rt_addr ? reg_26_3 : _GEN_153; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_155 = 5'h1b == io_Rt_addr ? reg_27_3 : _GEN_154; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_156 = 5'h1c == io_Rt_addr ? reg_28_3 : _GEN_155; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_157 = 5'h1d == io_Rt_addr ? reg_29_3 : _GEN_156; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_158 = 5'h1e == io_Rt_addr ? reg_30_3 : _GEN_157; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_159 = 5'h1f == io_Rt_addr ? reg_31_3 : _GEN_158; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_161 = 5'h1 == io_Rt_addr ? reg_1_2 : reg_0_2; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_162 = 5'h2 == io_Rt_addr ? reg_2_2 : _GEN_161; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_163 = 5'h3 == io_Rt_addr ? reg_3_2 : _GEN_162; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_164 = 5'h4 == io_Rt_addr ? reg_4_2 : _GEN_163; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_165 = 5'h5 == io_Rt_addr ? reg_5_2 : _GEN_164; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_166 = 5'h6 == io_Rt_addr ? reg_6_2 : _GEN_165; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_167 = 5'h7 == io_Rt_addr ? reg_7_2 : _GEN_166; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_168 = 5'h8 == io_Rt_addr ? reg_8_2 : _GEN_167; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_169 = 5'h9 == io_Rt_addr ? reg_9_2 : _GEN_168; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_170 = 5'ha == io_Rt_addr ? reg_10_2 : _GEN_169; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_171 = 5'hb == io_Rt_addr ? reg_11_2 : _GEN_170; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_172 = 5'hc == io_Rt_addr ? reg_12_2 : _GEN_171; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_173 = 5'hd == io_Rt_addr ? reg_13_2 : _GEN_172; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_174 = 5'he == io_Rt_addr ? reg_14_2 : _GEN_173; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_175 = 5'hf == io_Rt_addr ? reg_15_2 : _GEN_174; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_176 = 5'h10 == io_Rt_addr ? reg_16_2 : _GEN_175; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_177 = 5'h11 == io_Rt_addr ? reg_17_2 : _GEN_176; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_178 = 5'h12 == io_Rt_addr ? reg_18_2 : _GEN_177; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_179 = 5'h13 == io_Rt_addr ? reg_19_2 : _GEN_178; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_180 = 5'h14 == io_Rt_addr ? reg_20_2 : _GEN_179; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_181 = 5'h15 == io_Rt_addr ? reg_21_2 : _GEN_180; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_182 = 5'h16 == io_Rt_addr ? reg_22_2 : _GEN_181; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_183 = 5'h17 == io_Rt_addr ? reg_23_2 : _GEN_182; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_184 = 5'h18 == io_Rt_addr ? reg_24_2 : _GEN_183; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_185 = 5'h19 == io_Rt_addr ? reg_25_2 : _GEN_184; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_186 = 5'h1a == io_Rt_addr ? reg_26_2 : _GEN_185; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_187 = 5'h1b == io_Rt_addr ? reg_27_2 : _GEN_186; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_188 = 5'h1c == io_Rt_addr ? reg_28_2 : _GEN_187; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_189 = 5'h1d == io_Rt_addr ? reg_29_2 : _GEN_188; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_190 = 5'h1e == io_Rt_addr ? reg_30_2 : _GEN_189; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_191 = 5'h1f == io_Rt_addr ? reg_31_2 : _GEN_190; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_193 = 5'h1 == io_Rt_addr ? reg_1_1 : reg_0_1; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_194 = 5'h2 == io_Rt_addr ? reg_2_1 : _GEN_193; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_195 = 5'h3 == io_Rt_addr ? reg_3_1 : _GEN_194; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_196 = 5'h4 == io_Rt_addr ? reg_4_1 : _GEN_195; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_197 = 5'h5 == io_Rt_addr ? reg_5_1 : _GEN_196; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_198 = 5'h6 == io_Rt_addr ? reg_6_1 : _GEN_197; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_199 = 5'h7 == io_Rt_addr ? reg_7_1 : _GEN_198; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_200 = 5'h8 == io_Rt_addr ? reg_8_1 : _GEN_199; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_201 = 5'h9 == io_Rt_addr ? reg_9_1 : _GEN_200; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_202 = 5'ha == io_Rt_addr ? reg_10_1 : _GEN_201; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_203 = 5'hb == io_Rt_addr ? reg_11_1 : _GEN_202; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_204 = 5'hc == io_Rt_addr ? reg_12_1 : _GEN_203; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_205 = 5'hd == io_Rt_addr ? reg_13_1 : _GEN_204; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_206 = 5'he == io_Rt_addr ? reg_14_1 : _GEN_205; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_207 = 5'hf == io_Rt_addr ? reg_15_1 : _GEN_206; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_208 = 5'h10 == io_Rt_addr ? reg_16_1 : _GEN_207; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_209 = 5'h11 == io_Rt_addr ? reg_17_1 : _GEN_208; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_210 = 5'h12 == io_Rt_addr ? reg_18_1 : _GEN_209; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_211 = 5'h13 == io_Rt_addr ? reg_19_1 : _GEN_210; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_212 = 5'h14 == io_Rt_addr ? reg_20_1 : _GEN_211; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_213 = 5'h15 == io_Rt_addr ? reg_21_1 : _GEN_212; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_214 = 5'h16 == io_Rt_addr ? reg_22_1 : _GEN_213; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_215 = 5'h17 == io_Rt_addr ? reg_23_1 : _GEN_214; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_216 = 5'h18 == io_Rt_addr ? reg_24_1 : _GEN_215; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_217 = 5'h19 == io_Rt_addr ? reg_25_1 : _GEN_216; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_218 = 5'h1a == io_Rt_addr ? reg_26_1 : _GEN_217; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_219 = 5'h1b == io_Rt_addr ? reg_27_1 : _GEN_218; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_220 = 5'h1c == io_Rt_addr ? reg_28_1 : _GEN_219; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_221 = 5'h1d == io_Rt_addr ? reg_29_1 : _GEN_220; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_222 = 5'h1e == io_Rt_addr ? reg_30_1 : _GEN_221; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_223 = 5'h1f == io_Rt_addr ? reg_31_1 : _GEN_222; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [23:0] io_Rt_out_hi_1 = {_GEN_159,_GEN_191,_GEN_223}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_225 = 5'h1 == io_Rt_addr ? reg_1_0 : reg_0_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_226 = 5'h2 == io_Rt_addr ? reg_2_0 : _GEN_225; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_227 = 5'h3 == io_Rt_addr ? reg_3_0 : _GEN_226; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_228 = 5'h4 == io_Rt_addr ? reg_4_0 : _GEN_227; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_229 = 5'h5 == io_Rt_addr ? reg_5_0 : _GEN_228; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_230 = 5'h6 == io_Rt_addr ? reg_6_0 : _GEN_229; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_231 = 5'h7 == io_Rt_addr ? reg_7_0 : _GEN_230; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_232 = 5'h8 == io_Rt_addr ? reg_8_0 : _GEN_231; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_233 = 5'h9 == io_Rt_addr ? reg_9_0 : _GEN_232; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_234 = 5'ha == io_Rt_addr ? reg_10_0 : _GEN_233; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_235 = 5'hb == io_Rt_addr ? reg_11_0 : _GEN_234; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_236 = 5'hc == io_Rt_addr ? reg_12_0 : _GEN_235; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_237 = 5'hd == io_Rt_addr ? reg_13_0 : _GEN_236; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_238 = 5'he == io_Rt_addr ? reg_14_0 : _GEN_237; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_239 = 5'hf == io_Rt_addr ? reg_15_0 : _GEN_238; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_240 = 5'h10 == io_Rt_addr ? reg_16_0 : _GEN_239; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_241 = 5'h11 == io_Rt_addr ? reg_17_0 : _GEN_240; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_242 = 5'h12 == io_Rt_addr ? reg_18_0 : _GEN_241; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_243 = 5'h13 == io_Rt_addr ? reg_19_0 : _GEN_242; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_244 = 5'h14 == io_Rt_addr ? reg_20_0 : _GEN_243; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_245 = 5'h15 == io_Rt_addr ? reg_21_0 : _GEN_244; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_246 = 5'h16 == io_Rt_addr ? reg_22_0 : _GEN_245; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_247 = 5'h17 == io_Rt_addr ? reg_23_0 : _GEN_246; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_248 = 5'h18 == io_Rt_addr ? reg_24_0 : _GEN_247; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_249 = 5'h19 == io_Rt_addr ? reg_25_0 : _GEN_248; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_250 = 5'h1a == io_Rt_addr ? reg_26_0 : _GEN_249; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_251 = 5'h1b == io_Rt_addr ? reg_27_0 : _GEN_250; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_252 = 5'h1c == io_Rt_addr ? reg_28_0 : _GEN_251; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_253 = 5'h1d == io_Rt_addr ? reg_29_0 : _GEN_252; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_254 = 5'h1e == io_Rt_addr ? reg_30_0 : _GEN_253; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_255 = 5'h1f == io_Rt_addr ? reg_31_0 : _GEN_254; // @[Cat.scala 30:58 Cat.scala 30:58]
  assign io_Rs_out = {io_Rs_out_hi_1,_GEN_127}; // @[Cat.scala 30:58]
  assign io_Rt_out = {io_Rt_out_hi_1,_GEN_255}; // @[Cat.scala 30:58]
  always @(posedge clock) begin
    if (reset) begin // @[Register.scala 17:22]
      reg_0_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h0 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_0_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_0_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h0 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_0_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_0_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h0 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_0_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_0_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h0 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_0_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_1_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h1 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_1_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_1_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h1 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_1_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_1_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h1 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_1_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_1_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h1 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_1_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_2_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h2 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_2_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_2_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h2 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_2_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_2_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h2 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_2_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_2_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h2 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_2_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_3_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h3 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_3_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_3_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h3 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_3_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_3_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h3 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_3_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_3_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h3 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_3_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_4_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h4 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_4_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_4_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h4 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_4_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_4_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h4 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_4_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_4_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h4 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_4_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_5_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h5 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_5_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_5_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h5 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_5_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_5_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h5 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_5_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_5_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h5 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_5_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_6_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h6 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_6_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_6_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h6 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_6_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_6_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h6 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_6_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_6_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h6 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_6_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_7_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h7 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_7_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_7_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h7 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_7_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_7_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h7 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_7_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_7_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h7 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_7_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_8_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h8 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_8_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_8_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h8 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_8_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_8_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h8 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_8_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_8_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h8 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_8_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_9_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h9 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_9_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_9_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h9 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_9_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_9_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h9 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_9_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_9_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h9 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_9_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_10_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'ha == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_10_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_10_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'ha == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_10_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_10_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'ha == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_10_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_10_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'ha == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_10_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_11_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'hb == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_11_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_11_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'hb == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_11_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_11_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'hb == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_11_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_11_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'hb == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_11_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_12_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'hc == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_12_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_12_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'hc == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_12_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_12_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'hc == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_12_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_12_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'hc == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_12_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_13_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'hd == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_13_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_13_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'hd == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_13_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_13_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'hd == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_13_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_13_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'hd == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_13_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_14_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'he == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_14_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_14_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'he == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_14_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_14_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'he == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_14_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_14_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'he == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_14_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_15_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'hf == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_15_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_15_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'hf == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_15_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_15_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'hf == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_15_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_15_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'hf == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_15_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_16_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h10 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_16_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_16_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h10 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_16_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_16_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h10 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_16_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_16_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h10 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_16_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_17_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h11 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_17_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_17_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h11 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_17_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_17_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h11 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_17_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_17_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h11 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_17_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_18_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h12 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_18_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_18_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h12 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_18_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_18_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h12 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_18_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_18_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h12 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_18_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_19_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h13 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_19_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_19_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h13 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_19_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_19_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h13 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_19_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_19_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h13 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_19_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_20_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h14 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_20_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_20_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h14 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_20_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_20_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h14 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_20_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_20_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h14 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_20_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_21_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h15 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_21_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_21_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h15 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_21_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_21_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h15 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_21_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_21_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h15 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_21_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_22_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h16 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_22_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_22_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h16 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_22_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_22_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h16 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_22_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_22_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h16 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_22_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_23_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h17 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_23_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_23_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h17 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_23_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_23_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h17 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_23_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_23_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h17 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_23_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_24_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h18 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_24_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_24_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h18 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_24_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_24_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h18 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_24_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_24_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h18 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_24_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_25_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h19 == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_25_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_25_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h19 == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_25_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_25_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h19 == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_25_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_25_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h19 == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_25_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_26_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h1a == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_26_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_26_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h1a == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_26_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_26_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h1a == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_26_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_26_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h1a == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_26_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_27_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h1b == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_27_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_27_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h1b == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_27_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_27_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h1b == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_27_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_27_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h1b == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_27_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_28_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h1c == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_28_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_28_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h1c == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_28_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_28_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h1c == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_28_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_28_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h1c == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_28_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_29_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h1d == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_29_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_29_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h1d == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_29_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_29_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h1d == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_29_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_29_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h1d == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_29_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_30_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h1e == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_30_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_30_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h1e == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_30_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_30_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h1e == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_30_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_30_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h1e == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_30_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_31_0 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[0]) begin // @[Register.scala 22:33]
        if (5'h1f == io_Rd_addr) begin // @[Register.scala 23:32]
          reg_31_0 <= io_Rd_in[7:0]; // @[Register.scala 23:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_31_1 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[1]) begin // @[Register.scala 25:33]
        if (5'h1f == io_Rd_addr) begin // @[Register.scala 26:32]
          reg_31_1 <= io_Rd_in[15:8]; // @[Register.scala 26:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_31_2 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[2]) begin // @[Register.scala 28:33]
        if (5'h1f == io_Rd_addr) begin // @[Register.scala 29:32]
          reg_31_2 <= io_Rd_in[23:16]; // @[Register.scala 29:32]
        end
      end
    end
    if (reset) begin // @[Register.scala 17:22]
      reg_31_3 <= 8'h0; // @[Register.scala 17:22]
    end else if (io_Rd_addr != 5'h0) begin // @[Register.scala 21:29]
      if (io_Rd_byte_w_en[3]) begin // @[Register.scala 31:33]
        if (5'h1f == io_Rd_addr) begin // @[Register.scala 32:32]
          reg_31_3 <= io_Rd_in[31:24]; // @[Register.scala 32:32]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  reg_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  reg_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  reg_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  reg_1_0 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  reg_1_1 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  reg_1_2 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  reg_1_3 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  reg_2_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  reg_2_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  reg_2_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  reg_2_3 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  reg_3_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  reg_3_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  reg_3_2 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  reg_3_3 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  reg_4_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  reg_4_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  reg_4_2 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  reg_4_3 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  reg_5_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  reg_5_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  reg_5_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  reg_5_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  reg_6_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  reg_6_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  reg_6_2 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  reg_6_3 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  reg_7_0 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  reg_7_1 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  reg_7_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  reg_7_3 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  reg_8_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  reg_8_1 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  reg_8_2 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  reg_8_3 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  reg_9_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  reg_9_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  reg_9_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  reg_9_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  reg_10_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  reg_10_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  reg_10_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  reg_10_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  reg_11_0 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  reg_11_1 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  reg_11_2 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  reg_11_3 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  reg_12_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  reg_12_1 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  reg_12_2 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  reg_12_3 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  reg_13_0 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  reg_13_1 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  reg_13_2 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  reg_13_3 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  reg_14_0 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  reg_14_1 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  reg_14_2 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  reg_14_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  reg_15_0 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  reg_15_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  reg_15_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  reg_15_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  reg_16_0 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  reg_16_1 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  reg_16_2 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  reg_16_3 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  reg_17_0 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  reg_17_1 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  reg_17_2 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  reg_17_3 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  reg_18_0 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  reg_18_1 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  reg_18_2 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  reg_18_3 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  reg_19_0 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  reg_19_1 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  reg_19_2 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  reg_19_3 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  reg_20_0 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  reg_20_1 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  reg_20_2 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  reg_20_3 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  reg_21_0 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  reg_21_1 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  reg_21_2 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  reg_21_3 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  reg_22_0 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  reg_22_1 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  reg_22_2 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  reg_22_3 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  reg_23_0 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  reg_23_1 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  reg_23_2 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  reg_23_3 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  reg_24_0 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  reg_24_1 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  reg_24_2 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  reg_24_3 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  reg_25_0 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  reg_25_1 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  reg_25_2 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  reg_25_3 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  reg_26_0 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  reg_26_1 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  reg_26_2 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  reg_26_3 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  reg_27_0 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  reg_27_1 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  reg_27_2 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  reg_27_3 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  reg_28_0 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  reg_28_1 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  reg_28_2 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  reg_28_3 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  reg_29_0 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  reg_29_1 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  reg_29_2 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  reg_29_3 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  reg_30_0 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  reg_30_1 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  reg_30_2 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  reg_30_3 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  reg_31_0 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  reg_31_1 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  reg_31_2 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  reg_31_3 = _RAND_127[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
